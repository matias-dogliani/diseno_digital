 

/*La particion de un diseno digital en modulos es importante */

module top (
    
     input clock, 
     input i_reset, 
     input [3:0] i_sw,
     output [3:0] o_led,
     output [3:0] o_led_b,
     output [3:0] o_led_g
 
 );


 endmodule  




module top 
(
	
);

endmodule //top